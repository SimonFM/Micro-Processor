-- Simon Markham 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
entity control_memory_256 is
	port( MW, MM, RW, MD, MB, IL : out STD_LOGIC;
			TB, TA, TD, PL, PI, MC : out STD_LOGIC;
			FS : out STD_LOGIC_VECTOR(4 downto 0);
			MS : out STD_LOGIC_VECTOR(2 downto 0);
			NA : out STD_LOGIC_VECTOR(7 downto 0);
			IN_CAR : in STD_LOGIC_VECTOR(7 downto 0));
end control_memory_256;
architecture Behavioral of control_memory_256 is
	signal MWs, MMs, RWs, MDs, MBs, ILs : STD_LOGIC;
	signal TBs, TAs, TDs, PLs, PIs, MCs : STD_LOGIC;
	signal FSs : STD_LOGIC_VECTOR(4 downto 0);
	signal MSs : STD_LOGIC_VECTOR(2 downto 0);
	signal NAs : STD_LOGIC_VECTOR(7 downto 0);
	type mem_array is array(0 to 255) of STD_LOGIC_VECTOR(27 downto 0);
	begin
			memory_m: process(IN_CAR) 
			variable control_mem : mem_array:=(
													-- 0
													X"0018024", -- Messing around here
													X"0200024", -- ADD
													X"0200164", -- NOT
													X"0200014", -- INC
													X"0200001", -- ST
													X"020000C", -- LD
													X"0200144", -- ADI
													X"0300000", -- EXO
													X"000C002", -- IF
													X"0000009", -- 9
													X"000000A", -- A
													X"000000B", -- B
													X"000000C", -- C
													X"000000D", -- D
													X"000000E", -- E
													X"000000F", -- F
													-- 1
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 2
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 3
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 4
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 5
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 6
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 7
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 8
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 9
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 10
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 11
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 12
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 13
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 14
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000", -- F
													-- 14
													X"0000000", -- 0
													X"0000000", -- 1
													X"0000000", -- 2
													X"0000000", -- 3
													X"0000000", -- 4
													X"0000000", -- 5
													X"0000000", -- 6
													X"0000000", -- 7
													X"0000000", -- 8
													X"0000000", -- 9
													X"0000000", -- A
													X"0000000", -- B
													X"0000000", -- C
													X"0000000", -- D
													X"0000000", -- E
													X"0000000"); -- F	
			variable addr : integer;
			variable control_out : STD_LOGIC_VECTOR(27 downto 0);
			begin
					addr := CONV_INTEGER(IN_CAR);
					control_out := control_mem(addr);
					MW <= control_out(0);
					MM <= control_out(1);
					RW <= control_out(2);
					MD <= control_out(3);
					FS <= control_out(8 downto 4);
					MB <= control_out(9);
					TB <= control_out(10);
					TA <= control_out(11);
					TD <= control_out(12);
					PL <= control_out(13);
					PI <= control_out(14);
					IL <= control_out(15);
					MC <= control_out(16);
					MS <= control_out(19 downto 17);
					NA <= control_out(27 downto 20);
		  end process; 
end Behavioral;
